module riscv #(parameter width = 32,addrWidth = 5) (
	input clock,
	input	regWriteEnable,
	input	[addrWidth-1:0]addrA,
	input	[addrWidth-1:0]addrB,
	input [addrWidth-1:0]addrD,
	input [width-1:0]dataD,
	output [width-1:0]dataA,
	output [width-1:0]dataB
);
regFile rf(~clock,regWriteEnable,addrA,addrB,addrD,dataD,dataA,dataB);
endmodule








